// clock.v

// Generated using ACDS version 12.1 177 at 2022.07.22.10:15:19

`timescale 1 ps / 1 ps
module clock (
		output wire  clk_0_clk_clk,    //    clk_0_clk.clk
		input  wire  clk_0_clk_in_clk, // clk_0_clk_in.clk
		input  wire  reset_reset_n     //        reset.reset_n
	);

	assign clk_0_clk_clk = clk_0_clk_in_clk;

endmodule
