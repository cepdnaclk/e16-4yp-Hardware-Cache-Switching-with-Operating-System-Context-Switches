module instruction_decode_unit (
   
);
    
endmodule