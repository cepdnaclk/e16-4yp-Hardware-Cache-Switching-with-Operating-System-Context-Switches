// pll.v

// Generated using ACDS version 12.1 177 at 2022.07.22.10:20:40

`timescale 1 ps / 1 ps
module pll (
		input  wire  reset_1_reset,    //      reset_1.reset
		output wire  clock_output_clk, // clock_output.clk
		input  wire  clock_input_clk   //  clock_input.clk
	);

	pll_altpll_0 altpll_0 (
		.clk       (clock_input_clk),  //       inclk_interface.clk
		.reset     (reset_1_reset),    // inclk_interface_reset.reset
		.read      (),                 //             pll_slave.read
		.write     (),                 //                      .write
		.address   (),                 //                      .address
		.readdata  (),                 //                      .readdata
		.writedata (),                 //                      .writedata
		.c0        (clock_output_clk), //                    c0.clk
		.areset    (),                 //        areset_conduit.export
		.locked    (),                 //        locked_conduit.export
		.phasedone ()                  //     phasedone_conduit.export
	);

endmodule
